netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float EntMM29lc_lai_for_1kmx1km(lat, lon) ;
		EntMM29lc_lai_for_1kmx1km:long_name = "EntMM 29 lc_lai_for_1kmx1km check sum cover" ;
}
