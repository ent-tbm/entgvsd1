netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float drought_br(lat, lon) ;
		drought_br:long_name = "7 - drought deciduous broadleaf EntMM LAI max 1kmx1km" ;
}
