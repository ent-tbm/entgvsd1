netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float crops_c3_herb(lat, lon) ;
		crops_c3_herb:long_name = "15 - crops C3 herb EntMM LAI max 1kmx1km" ;
}
