netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float decid_nd(lat, lon) ;
		decid_nd:long_name = "8 - deciduous needleleaf EntMM LAI max 1kmx1km" ;
}
