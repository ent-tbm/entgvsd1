netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float EntdominantPFT_check_sum_Jun_1kmx1km(lat, lon) ;
		EntdominantPFT_check_sum_Jun_1kmx1km:long_name = "Ent dominant PFT check sum Jun 1kmx1km" ;
}
