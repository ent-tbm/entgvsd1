netcdf EntPFTs_percell_check_sum_Jun_1kmx1km {
dimensions:
        lon = 43200 ;
        lat = 21600 ;

variables:
        float lon(lon) ;
        float lat(lat) ;

        float EntPFTs_percell_check_sum_Jun_1kmx1km(lat, lon) ;
            EntPFTs_percell_check_sum_Jun_1kmx1km:long_name = "Ent PFTs per cell check sum Jun 1kmx1km" ;

}

