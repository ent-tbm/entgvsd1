netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float water_lc(lat, lon) ;
		water_lc:long_name = "WATER (cover fraction)" ;
}
