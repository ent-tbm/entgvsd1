netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float ever_br_late(lat, lon) ;
		ever_br_late:long_name = "2 - evergreen broadleaf late successional" ;
}
