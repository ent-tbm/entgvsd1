netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float bare_sparse(lat, lon) ;
		bare_sparse:long_name = "19 - Bare or sparsely vegetated, urban" ;
}
