netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float ever_nd_late(lat, lon) ;
		ever_nd_late:long_name = "4 - evergreen needleleaf late successional" ;
}
