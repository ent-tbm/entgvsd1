netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float ever_br_early(lat, lon) ;
		ever_br_early:long_name = "1 - evergreen broadleaf early successional EntMM LAI max 1kmx1km" ;
}
