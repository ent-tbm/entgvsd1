netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float c3_grass_ann(lat, lon) ;
		c3_grass_ann:long_name = "13 - C3 grass - annual EntMM LAI max 1kmx1km" ;
}
