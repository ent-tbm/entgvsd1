netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float crops_c4_herb(lat, lon) ;
		crops_c4_herb:long_name = "16 - crops C4 herb EntMM LAI max 1kmx1km" ;
}
