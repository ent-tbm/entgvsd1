netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float lon(lon) ;
	float lat(lat) ;
	float snow_ice(lat, lon) ;
		snow_ice:long_name = "18 - Permanent snow/ice" ;
}
