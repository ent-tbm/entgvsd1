netcdf x {
dimensions:
	lon = 43200 ;
	lat = 21600 ;
variables:
	float EntLAI_check_sum_Jun_1kmx1km(lat, lon) ;
		EntLAI_check_sum_Jun_1kmx1km:long_name = "Ent LAI check sum Jun 1kmx1km" ;
}
